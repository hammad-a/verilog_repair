/////////////////////////////////////////////////////////////////////////
//                                                                     //
//   Modulename :  sys_defs.vh                                         //
//                                                                     //
//  Description :  This file has the parameter and typedefs used in    //
//                 in-lab 3 part b                                     //
//                                                                     //
/////////////////////////////////////////////////////////////////////////

typedef enum {WAIT, WATCH, ASSERT} STATE;
typedef enum {RAND, MATCH, NO_MATCH} OVERRIDE;

parameter CLOCK_PERIOD = 10;
